library ieee;
use ieee.std_logic_1164.all;

entity control is
	ctrl1, ctrl2, ctrl3: in std_logic;
end entity;

architecture bhvr of control is

	signal -- completar

begin
end architecture;