library ieee;
use ieee.std_logic_1164.all;

entity leituraRAM is

end entity;

architecture bhvr of leituraRAM is
begin
end architecture;