-- apenas vamos declarar e usar o arquivo 
-- presente no moodle