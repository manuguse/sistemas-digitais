library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity registerN is
	generic(	width: natural;
				resetValue: integer := 0 );
	port(	-- control
			clock, reset, load: in std_logic;
			-- data
			input: in std_logic_vector(width-1 downto 0);
			output: out std_logic_vector(width-1 downto 0));
end entity;

architecture behav0 of registerN is
    signal currentState, nextState: std_logic_vector(width-1 downto 0);
begin
    -- next-state logic  (nao exclua e nem mude esta linha)
    nextState <= input when load = '1' else currentState;

	-- memory element --state register-- (nao exclua e nem mude esta linha)
    process(clock, reset)
    begin
        if reset = '1' then
            output <= std_logic_vector(to_unsigned(resetValue, width));
        elsif rising_edge(clock) then
            if load = '1' then
                currentState <= nextState;
            end if;
        end if;
    end process;
	
	-- output logic  (nao exclua e nem mude esta linha)
	output <= currentState;
end architecture;