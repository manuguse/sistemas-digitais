library ieee;
use ieee.std_logic_1164.all;

entity datapath is
port();

end entity;

architecture bhvr of datapath is

	signal -- completar

begin
end architecture;